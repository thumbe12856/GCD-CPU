`define IM_MAX 256
`define IMSIZE 8
`timescale 1ns/1ps

module INSTRUCTION_MEMORY(
	clk,
	wea,
	addr,
	din,
	dout
);

input clk, wea;
input [`IMSIZE-1:0] addr;
input [31:0] din;

output [31:0] dout;

// IM_MAX = how many memory space can use
reg [31:0] instruction [0:`IM_MAX-1];

initial
begin

	instruction[0] = 32'b000000_00000_00000_00000_00000_100000;		//NOP(add $0, $0, $0)
	instruction[1] = 32'b000000_00000_00000_00000_00000_100000;		//NOP(add $0, $0, $0)

	//lw $t1, 0($0)
	instruction[2] = 32'b100011_00000_01001_00000_00000_000000;		//lw $9, 0($0) , first num

	//lw $t2, 4($0)
	instruction[3] = 32'b100011_00000_01010_00000_00000_000100;		//lw $10, 4($0) , second num
	instruction[4] = 32'b000000_00000_00000_00000_00000_100010;		//NOP(sub $0, $0, $0)
	instruction[5] = 32'b000000_00000_00000_00000_00000_100000;		//NOP(add $0, $0, $0)
	instruction[6] = 32'b000000_00000_00000_00000_00000_100000;		//NOP(add $0, $0, $0)

	//GCD
	//sub $sp, $sp, 4
	instruction[7] = 32'b000000_11101_00010_11101_00000_100010; 	//sub $29, $29, $2
	instruction[8] = 32'b000000_00000_00000_00000_00000_100010; 	//NOP(sub $0, $0, $0)
	instruction[9] = 32'b000000_00000_00000_00000_00000_100000;		//NOP(add $0, $0, $0)
	instruction[10] = 32'b000000_00000_00000_00000_00000_100000; 	//NOP(add $0, $0, $0)

	//sw $ra, 0($sp)
	instruction[11] = 32'b101011_11101_11111_00000_00000_000000; 	//sw $31, 0($29)
	instruction[12] = 32'b000000_00000_00000_00000_00000_100010; 	//NOP(sub $0, $0, $0)
	instruction[13] = 32'b000000_00000_00000_00000_00000_100000; 	//NOP(add $0, $0, $0)
	instruction[14] = 32'b000000_00000_00000_00000_00000_100000; 	//NOP(add $0, $0, $0)

	//beq $t1, $t2, GCD_is_t1:34
	instruction[15] = 32'b000100_01001_01010_00000_00000_010010;	//beq $9 $10 18
	instruction[16] = 32'b000000_00000_00000_00000_00000_100010;	//NOP(sub $0, $0, $0)
	instruction[17] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	instruction[18] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	instruction[19] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)

	//beq $t1, $t3, GCD_is_one:42
	instruction[20] = 32'b000100_01001_00001_00000_00000_010101;	//beq $9 $1 21
	instruction[21] = 32'b000000_00000_00000_00000_00000_100010;	//NOP(sub $0, $0, $0)
	instruction[22] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	instruction[23] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	instruction[24] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)

	//beq $t2, $t3, GCD_is_one:42
	instruction[25] = 32'b000100_01010_00001_00000_00000_010000;	//beq $10 $1 16
	instruction[26] = 32'b000000_00000_00000_00000_00000_100010;	//NOP(sub $0, $0, $0)
	instruction[27] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	instruction[28] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	instruction[29] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)

	//j Deal_number:50
	instruction[30] = 32'b000010_00000_00000_00000_00000_110010; 	//j 50
	instruction[31] = 32'b000000_00000_00000_00000_00000_100010;	//NOP(sub $0, $0, $0)
	instruction[32] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	instruction[33] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)

	//GCD_is_t1
	//sw $t1, 8($zero)
	instruction[34] = 32'b101011_00000_01001_00000_00000_001000; 	//sw $9, 8($0)
	//instruction[35] = 32'b000000_00000_00000_00000_00000_100010; 	//NOP(sub $0, $0, $0)
	instruction[35] = 32'b000000_00000_00000_00000_00000_100010;	//NOP(sub $0, $0, $0)
	instruction[36] = 32'b000000_00000_00000_00000_00000_100000; 	//NOP(add $0, $0, $0)
	instruction[37] = 32'b000000_00000_00000_00000_00000_100000; 	//NOP(add $0, $0, $0)

	//jr $ra
	instruction[38] = 32'b000000_11111_00000_00000_00000_001000; 	//jr r31
	instruction[39] = 32'b000000_00000_00000_00000_00000_100010; 	//NOP(sub $0, $0, $0)
	instruction[40] = 32'b000000_00000_00000_00000_00000_100000; 	//NOP(add $0, $0, $0)
	instruction[41] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)

	//GCD_is_one
	//sw $t3, 8($zero)
	instruction[42] = 32'b101011_00000_00001_00000_00000_001000; 	//sw $1, 8($0)
	instruction[43] = 32'b000000_00000_00000_00000_00000_100010; 	//NOP(sub $0, $0, $0)
	instruction[44] = 32'b000000_00000_00000_00000_00000_100000; 	//NOP(add $0, $0, $0)
	instruction[45] = 32'b000000_00000_00000_00000_00000_100000; 	//NOP(add $0, $0, $0)

	//jr $ra
	instruction[46] = 32'b000000_11111_00000_00000_00000_001000; 	//jr r31
	instruction[47] = 32'b000000_00000_00000_00000_00000_100010; 	//NOP(sub $0, $0, $0)
	instruction[48] = 32'b000000_00000_00000_00000_00000_100000; 	//NOP(add $0, $0, $0)
	instruction[49] = 32'b000000_00000_00000_00000_00000_100000; 	//NOP(add $0, $0, $0)

	//Deal_number
	//slt $t0, $t1, $t2	-> t1 < t2 ? 1 : 0
	instruction[50] = 32'b000000_01001_01010_01000_00000_101010;	//slt $8, $9, $10 :  $8 = $9 < $10 ? 1 : 0
	instruction[51] = 32'b000000_00000_00000_00000_00000_100010;	//NOP(sub $0, $0, $0)
	instruction[52] = 32'b000000_00000_00000_00000_00000_100010;	//NOP(sub $0, $0, $0)
	instruction[53] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	instruction[54] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)

	//beq $t0, $t3, t2_is_big:72
	instruction[55] = 32'b000100_01000_00001_00000_00000_010000;	//beq $8 $1 16
	instruction[56] = 32'b000000_00000_00000_00000_00000_100010;	//NOP(sub $0, $0, $0)
	instruction[57] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	instruction[58] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	instruction[59] = 32'b000000_00000_00000_00000_00000_100000;		//NOP(add $0, $0, $0)


	//t1_is_big
	//sub $t1, $t1, $t2
	instruction[60] = 32'b000000_01001_01010_01001_00000_100010;	//sub $9, $9, $10
	instruction[61] = 32'b000000_00000_00000_00000_00000_100010;	//NOP(sub $0, $0, $0)
	instruction[62] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	instruction[63] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)

	//jal GCD:7
	instruction[64] = 32'b000011_00000_00000_00000_00000_000111; 	//jal 7
	instruction[65] = 32'b000000_00000_00000_00000_00000_100000; 	//NOP(add $0, $0, $0)
	instruction[66] = 32'b000000_00000_00000_00000_00000_100000; 	//NOP(add $0, $0, $0)
	instruction[67] = 32'b000000_00000_00000_00000_00000_100000; 	//NOP(add $0, $0, $0)

	//j print_data:80
	instruction[68] = 32'b000010_00000_00000_00000_00001_010000; 	//j 80
	instruction[69] = 32'b000000_00000_00000_00000_00000_100010;	//NOP(sub $0, $0, $0)
	instruction[70] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	instruction[71] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)

	//t2_is_big
	//sub $t2, $t2, $t1
	instruction[72] = 32'b000000_01010_01001_01010_00000_100010;	//sub $10, $10, $9
	instruction[73] = 32'b000000_00000_00000_00000_00000_100010;	//NOP(sub $0, $0, $0)
	instruction[74] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	instruction[75] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)

	//jal GCD:7
	instruction[76] = 32'b000011_00000_00000_00000_00000_000111; 	//jal 7
	instruction[77] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	instruction[78] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	instruction[79] = 32'b000000_00000_00000_00000_00000_100000; 	//NOP(add $0, $0, $0)

	//print_data
	//lw $ra, 0($sp)
	instruction[80] = 32'b100011_11101_11111_00000_00000_000000;	//lw $31, 0($29)

	//addi $sp,$sp,4
	instruction[81] = 32'b000000_11101_00100_11101_00000_100000;	//add $29, $29, $4
	instruction[82] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	instruction[83] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	instruction[84] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)

	//jr $ra
	instruction[85] = 32'b000000_11111_00000_00000_00000_001000; 	//jr r31
	instruction[86] = 32'b000000_00000_00000_00000_00000_100010; 	//NOP(sub $0, $0, $0)
	instruction[87] = 32'b000000_00000_00000_00000_00000_100000; 	//NOP(add $0, $0, $0)
	instruction[88] = 32'b000000_00000_00000_00000_00000_100000; 	//NOP(add $0, $0, $0)
	
end



reg [`IMSIZE-1:0] addr_reg;

// if memory can use, then direct output
assign dout = instruction[addr_reg] ;

// for outside write instruction
always @(posedge clk)
begin
	//$display("------IM: dout:%b", dout);
	addr_reg <= addr[`IMSIZE-1:0];
	if(wea)
		instruction[addr[`IMSIZE-1:0]] <= din;
end

endmodule

